module reg_file(

);
    
endmodule