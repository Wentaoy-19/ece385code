module ALU(
    
);
    
endmodule