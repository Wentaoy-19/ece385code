module datapath(
input logic Clk,
input logic Reset_ah, Continue_ah, Run_ah, 
input logic BEN,LD_MAR,LD_MDR,LD_IR,LD_BEN,LD_CC,LD_REG,LD_PC,LD_LED,
input logic GatePC, GateMDR, GateALU,GateMARMUX,
input logic[1:0] PCMUX,ADDR2MUX,ALUK,
input logic DRMUX, SR1MUX, SR2MUX, ADDR1MUX,
input logic MIO_EN,
input logic[15:0] MDR_In, MAR, MDR, IR, PC,Data_from_SRAM, Data_to_SRAM
); // TODO:input ? output? 

logic[15:0] BUS;

logic[15:0] MDR_input;

always_ff @(posedge Clk) begin

end



always_comb begin
    if(MIO_EN)

end

endmodule